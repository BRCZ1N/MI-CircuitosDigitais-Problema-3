//------------------------------------------------------------------------------
//	Module:		LevelToPulseMealy
//	Desc:		This module provides a 1-cycle output based on a push button
//				raw input source.
//	Params:		This module is not parameterized.
//	Inputs:		See Lab2 document
//	Outputs:	See Lab2 document
//
//	Author:     YOUR NAME GOES HERE
//------------------------------------------------------------------------------
module	LevelToPulseMealy(
			//------------------------------------------------------------------
			//	Clock & Reset Inputs
			//------------------------------------------------------------------
			Clock,
			Reset,
			//------------------------------------------------------------------
			
			//------------------------------------------------------------------
			//	Inputs
			//------------------------------------------------------------------
			Level,
			//------------------------------------------------------------------
			
			//------------------------------------------------------------------
			//	Outputs
			//------------------------------------------------------------------
			Pulse
			//------------------------------------------------------------------
	);
	//--------------------------------------------------------------------------
	//	Clock & Reset Inputs
	//--------------------------------------------------------------------------
	input					Clock;	// System clock
	input					Reset;	// System reset
	//--------------------------------------------------------------------------
	
	//--------------------------------------------------------------------------
	//	Inputs
	//--------------------------------------------------------------------------
	input					Level;
	//--------------------------------------------------------------------------

	//--------------------------------------------------------------------------
	//	Outputs
	//--------------------------------------------------------------------------
	output					Pulse;
	//--------------------------------------------------------------------------

	//--------------------------------------------------------------------------
	//	State Encoding
	//--------------------------------------------------------------------------
	
	
	//--------------------------------------------------------------------------
	//	Wire Declarations
	//--------------------------------------------------------------------------
	
	wire D;
	
	//--------------------------------------------------------------------------
	
	//-------------------------------------------------------------------------
	//	Logic
	//--------------------------------------------------------------------------

	assign D	= Level;
	
	modulo_divisor_frequencia(.clr(),.clk(Clock),.clk_div(clk_div_r));
	
	modulo_ff_d ff_1(.d(Level),.clk(clk_div_r),.clr(Reset),.q(Qi),.nq());
	
	not(NQi,Qi);
	
	and(Pulse,Level,NQi);
		

	//--------------------------------------------------------------------------
endmodule // LevelToPulseMealy