//------------------------------------------------------------------------------
//	Module:		LevelToPulse
//	Desc:		This module provides a 1-cycle output based on a push button
//				raw input source.
//	Params:		This module is not parameterized.
//	Inputs:		See Lab2 document
//	Outputs:	See Lab2 document
//
//	Author:     YOUR NAME GOES HERE
//------------------------------------------------------------------------------
module	LevelToPulseMoore(
			//------------------------------------------------------------------
			//	Clock & Reset Inputs
			//------------------------------------------------------------------
			Clock,
			Reset,
			//------------------------------------------------------------------
			
			//------------------------------------------------------------------
			//	Inputs
			//------------------------------------------------------------------
			Level,
			//------------------------------------------------------------------
			
			//------------------------------------------------------------------
			//	Outputs
			//------------------------------------------------------------------
			Pulse
			//------------------------------------------------------------------
	);
	//--------------------------------------------------------------------------
	//	Clock & Reset Inputs
	//--------------------------------------------------------------------------
	input					Clock;	// System clock
	input					Reset;	// System reset
	//--------------------------------------------------------------------------
	
	//--------------------------------------------------------------------------
	//	Inputs
	//--------------------------------------------------------------------------
	input					Level;
	//--------------------------------------------------------------------------

	//--------------------------------------------------------------------------
	//	Outputs
	//--------------------------------------------------------------------------
	output					Pulse;
	//--------------------------------------------------------------------------

	//--------------------------------------------------------------------------
	//	State Encoding
	//--------------------------------------------------------------------------
	
	// place state encoding here
	
	//--------------------------------------------------------------------------
	
	//--------------------------------------------------------------------------
	//	Wire Declarations
	//--------------------------------------------------------------------------
	
	wire D0;
	wire D1;
	wire clk_div_r;
	wire NQi1;
	
	//--------------------------------------------------------------------------
	
	//--------------------------------------------------------------------------
	//	Logic
	//--------------------------------------------------------------------------

	and(D1,Level,Qi0);
	assign D0 = Level;
	
	modulo_divisor_frequencia(.clr(),.clk(Clock),.clk_div(clk_div_r));
	
	modulo_ff_d ff_1(.d(D1),.clk(clk_div_r),.clr(Reset),.q(Qi1),.nq());
	
	modulo_ff_d ff_2(.d(Level),.clk(clk_div_r),.clr(Reset),.q(Qi0),.nq());
	
	not(NQi1,Qi1);
	
	and(Pulse,NQi1,Qi0);
	

	//--------------------------------------------------------------------------
endmodule // LevelToPulse